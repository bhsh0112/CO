`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:45:49 11/14/2023 
// Design Name: 
// Module Name:    E_jump 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module E_jump(
    input [15:0] E_imm16,
    input [25:0] E_imm26,
    output [31:0] E_imm16_EXT,
    output [31:0] E_imm26_EXT
    );


endmodule
